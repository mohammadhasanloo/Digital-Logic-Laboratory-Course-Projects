library verilog;
use verilog.vl_types.all;
entity PWM_TB is
end PWM_TB;
