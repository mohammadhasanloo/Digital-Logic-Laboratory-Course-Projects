library verilog;
use verilog.vl_types.all;
entity DDS_TB is
end DDS_TB;
