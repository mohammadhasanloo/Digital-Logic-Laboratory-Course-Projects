library verilog;
use verilog.vl_types.all;
entity Waveform_Generator_TB is
end Waveform_Generator_TB;
