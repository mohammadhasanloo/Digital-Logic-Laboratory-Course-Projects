library verilog;
use verilog.vl_types.all;
entity Amplitute_Selector_TB is
end Amplitute_Selector_TB;
