library verilog;
use verilog.vl_types.all;
entity Frequency_Selector_TB is
end Frequency_Selector_TB;
