module Amplitute_Selector(in, SW, out);
  input [7:0] in;
  input[1:0] SW;
  output reg [7:0] out;
  
  always@(in, SW) begin
    if(SW==2'b00)
      out <= in;
    else if(SW==2'b01)
      out <= in >>> 1;
    else if(SW==2'b10)
      out <= in >>> 2;   
    else if(SW==2'b11)
      out <= in >>> 3;  
  end
endmodule