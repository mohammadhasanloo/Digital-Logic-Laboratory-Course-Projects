module wrapper_counter #(parameter N = 5) (
    input clk, rst, inc,
    output reg [7:0] count,
    output co
);
    always @(posedge clk or posedge rst) begin
        
        if (rst) count <= 8'b0;
        else if (inc) begin
            if (co) count <= 8'b0;
            else count <= count + 8'b00000001;
        end
    end

    assign co = (count == N - 1);
endmodule
