`timescale 1ns/1ns

module Waveform_Generator (input clk , rst , input [2:0]func , input [7:0]count_num , output reg [7:0]waveform);
    
    
    reg [7:0] reciprocal , square , triangle , dds;
	wire [7:0] sine , full_wave_rectified , half_wave_rectified;
    reg [15:0] curr_sin , oldCos , curr_cos , oldSine;

    // SQUARE
    always @(posedge clk) begin
        if (rst)
            square = 0;
        else begin
            if (count_num[7])
              square = 255;   
            else
              square = 0;
        end
    end
    
    // TRIANGLE
    always @(posedge clk) begin
        if (rst)
            triangle = 0;
        else begin
            if (count_num[7])
                triangle = triangle - 1'b1;
            else
                triangle = triangle + 1'b1;
        end
    end
    
    // RECIPROCAL
    always @(posedge clk) begin
        if(rst)
            reciprocal = 0;
        else
            reciprocal = (255 / (255 - count_num));
    end

    // SINE
    always @(posedge clk, posedge rst) begin
        if(rst) begin
            oldCos <= 16'd30000;
            oldSine <= 16'd0;
        end
        else begin
            oldCos <= curr_cos;
            oldSine <= curr_sin;

        end
    end

    always @(oldSine, oldCos) begin
        curr_sin = oldSine + {{6{oldCos[15]}}, oldCos[15:6]};
        curr_cos = oldCos - {{6{curr_sin[15]}}, curr_sin[15:6]};

    end

    assign sine = curr_sin[15:8];
    
    // FILL_WAVED
    assign full_wave_rectified = curr_sin[15] == 1 ? ~curr_sin[15:8]+1 : curr_sin[15:8];
    // HALF_WAVED
    assign half_wave_rectified = curr_sin[15] == 1 ? 8'b0 : curr_sin[15:8];


    always @(posedge clk) begin
        case (func)
            3'b000 : waveform = reciprocal;
            3'b001 : waveform = square ;
            3'b010 : waveform = triangle ;
            3'b011 : waveform = sine ;
            3'b100 : waveform = full_wave_rectified ;
            3'b101 : waveform = half_wave_rectified ;
            3'b110 : waveform = dds ;
        endcase
    end
    
endmodule
    
