library verilog;
use verilog.vl_types.all;
entity wg_test is
end wg_test;
