library verilog;
use verilog.vl_types.all;
entity exponential_TB is
end exponential_TB;
