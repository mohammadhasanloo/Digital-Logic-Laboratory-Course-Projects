library verilog;
use verilog.vl_types.all;
entity wgp_test is
end wgp_test;
